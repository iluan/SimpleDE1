	library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

ENTITY overwrap IS
PORT(
---------FPGA Connections-------------
CLOCK_50: IN STD_LOGIC;
---------HPS Connections---------------
HPS_CONV_USB_N:INOUT STD_LOGIC;
HPS_DDR3_ADDR:OUT STD_LOGIC_VECTOR(14 downto 0);
HPS_DDR3_BA: OUT STD_LOGIC_VECTOR(2 downto 0);
HPS_DDR3_CAS_N: OUT STD_LOGIC;
HPS_DDR3_CKE:OUT STD_LOGIC;
HPS_DDR3_CK_N: OUT STD_LOGIC;
HPS_DDR3_CK_P: OUT STD_LOGIC;
HPS_DDR3_CS_N: OUT STD_LOGIC;
HPS_DDR3_DM: OUT STD_LOGIC_VECTOR(3 downto 0);
HPS_DDR3_DQ: INOUT STD_LOGIC_VECTOR(31 downto 0);
HPS_DDR3_DQS_N: INOUT STD_LOGIC_VECTOR(3 downto 0);
HPS_DDR3_DQS_P: INOUT STD_LOGIC_VECTOR(3 downto 0);
HPS_DDR3_ODT: OUT STD_LOGIC;
HPS_DDR3_RAS_N: OUT STD_LOGIC;
HPS_DDR3_RESET_N: OUT  STD_LOGIC;
HPS_DDR3_RZQ: IN  STD_LOGIC;
HPS_DDR3_WE_N: OUT STD_LOGIC;
HPS_ENET_GTX_CLK: OUT STD_LOGIC;
HPS_ENET_INT_N:INOUT STD_LOGIC;
HPS_ENET_MDC:OUT STD_LOGIC;
HPS_ENET_MDIO:INOUT STD_LOGIC;
HPS_ENET_RX_CLK: IN STD_LOGIC;
HPS_ENET_RX_DATA: IN STD_LOGIC_VECTOR(3 downto 0);
HPS_ENET_RX_DV: IN STD_LOGIC;
HPS_ENET_TX_DATA: OUT STD_LOGIC_VECTOR(3 downto 0);
HPS_ENET_TX_EN: OUT STD_LOGIC;
HPS_KEY: INOUT STD_LOGIC;
HPS_SD_CLK: OUT STD_LOGIC;
HPS_SD_CMD: INOUT STD_LOGIC;
HPS_SD_DATA: INOUT STD_LOGIC_VECTOR(3 downto 0);
HPS_UART_RX: IN   STD_LOGIC;
HPS_UART_TX: OUT STD_LOGIC;
HPS_USB_CLKOUT: IN STD_LOGIC;
HPS_USB_DATA:INOUT STD_LOGIC_VECTOR(7 downto 0);
HPS_USB_DIR: IN STD_LOGIC;
HPS_USB_NXT: IN STD_LOGIC;
HPS_USB_STP: OUT STD_LOGIC

);
END overwrap;

ARCHITECTURE MAIN OF Overwrap IS
component WRAP0 is
	port ( 
		--Copia aquí los puertos de Wrap0
	);
end component;


	 component SIMPLE IS
PORT(
---------FPGA Connections-------------
CLOCK_50: IN STD_LOGIC;
init:OUT STD_LOGIC_VECTOR(7 downto 0);
count: IN UNSIGNED(7 downto 0);
---------HPS Connections---------------
HPS_CONV_USB_N:INOUT STD_LOGIC;
HPS_DDR3_ADDR:OUT STD_LOGIC_VECTOR(14 downto 0);
HPS_DDR3_BA: OUT STD_LOGIC_VECTOR(2 downto 0);
HPS_DDR3_CAS_N: OUT STD_LOGIC;
HPS_DDR3_CKE:OUT STD_LOGIC;
HPS_DDR3_CK_N: OUT STD_LOGIC;
HPS_DDR3_CK_P: OUT STD_LOGIC;
HPS_DDR3_CS_N: OUT STD_LOGIC;
HPS_DDR3_DM: OUT STD_LOGIC_VECTOR(3 downto 0);
HPS_DDR3_DQ: INOUT STD_LOGIC_VECTOR(31 downto 0);
HPS_DDR3_DQS_N: INOUT STD_LOGIC_VECTOR(3 downto 0);
HPS_DDR3_DQS_P: INOUT STD_LOGIC_VECTOR(3 downto 0);
HPS_DDR3_ODT: OUT STD_LOGIC;
HPS_DDR3_RAS_N: OUT STD_LOGIC;
HPS_DDR3_RESET_N: OUT  STD_LOGIC;
HPS_DDR3_RZQ: IN  STD_LOGIC;
HPS_DDR3_WE_N: OUT STD_LOGIC;
HPS_ENET_GTX_CLK: OUT STD_LOGIC;
HPS_ENET_INT_N:INOUT STD_LOGIC;
HPS_ENET_MDC:OUT STD_LOGIC;
HPS_ENET_MDIO:INOUT STD_LOGIC;
HPS_ENET_RX_CLK: IN STD_LOGIC;
HPS_ENET_RX_DATA: IN STD_LOGIC_VECTOR(3 downto 0);
HPS_ENET_RX_DV: IN STD_LOGIC;
HPS_ENET_TX_DATA: OUT STD_LOGIC_VECTOR(3 downto 0);
HPS_ENET_TX_EN: OUT STD_LOGIC;
HPS_KEY: INOUT STD_LOGIC;
HPS_SD_CLK: OUT STD_LOGIC;
HPS_SD_CMD: INOUT STD_LOGIC;
HPS_SD_DATA: INOUT STD_LOGIC_VECTOR(3 downto 0);
HPS_UART_RX: IN   STD_LOGIC;
HPS_UART_TX: OUT STD_LOGIC;
HPS_USB_CLKOUT: IN STD_LOGIC;
HPS_USB_DATA:INOUT STD_LOGIC_VECTOR(7 downto 0);
HPS_USB_DIR: IN STD_LOGIC;
HPS_USB_NXT: IN STD_LOGIC;
HPS_USB_STP: OUT STD_LOGIC
);
end component simple;
SIGNAL HPS_H2F_RST:STD_LOGIC;
--inserta aquí las señales que conectan a tu componente
BEGIN
u0: component WRAP0
	port map(
		--inserta aquí el mapa de puertos de wrap
	);

--FROM_HPS(7 downto 6) <= 'x';
u1 : component simple
        port map (
				---------FPGA Connections-------------
--CLOCK_50	=>	CLOCK_50,
--Aquí pon cualquier conexión entre el FPGA y el HPS
---------HPS Connections---------------
HPS_CONV_USB_N	=>	HPS_CONV_USB_N,
HPS_DDR3_ADDR	=>	HPS_DDR3_ADDR,
HPS_DDR3_BA	=>	HPS_DDR3_BA,
HPS_DDR3_CAS_N	=>	HPS_DDR3_CAS_N,
HPS_DDR3_CKE	=>	HPS_DDR3_CKE,
HPS_DDR3_CK_N	=>	HPS_DDR3_CK_N,
HPS_DDR3_CK_P	=>	HPS_DDR3_CK_P,
HPS_DDR3_CS_N	=>	HPS_DDR3_CS_N,
HPS_DDR3_DM	=>	HPS_DDR3_DM,
HPS_DDR3_DQ	=>	HPS_DDR3_DQ,
HPS_DDR3_DQS_N	=>	HPS_DDR3_DQS_N,
HPS_DDR3_DQS_P	=>	HPS_DDR3_DQS_P,
HPS_DDR3_ODT	=>	HPS_DDR3_ODT,
HPS_DDR3_RAS_N	=>	HPS_DDR3_RAS_N,
HPS_DDR3_RESET_N	=>	HPS_DDR3_RESET_N,
HPS_DDR3_RZQ	=>	HPS_DDR3_RZQ,
HPS_DDR3_WE_N	=>	HPS_DDR3_WE_N,
HPS_ENET_GTX_CLK	=>	HPS_ENET_GTX_CLK,
HPS_ENET_INT_N	=>	HPS_ENET_INT_N,
HPS_ENET_MDC	=>	HPS_ENET_MDC,
HPS_ENET_MDIO	=>	HPS_ENET_MDIO,
HPS_ENET_RX_CLK	=>	HPS_ENET_RX_CLK,
HPS_ENET_RX_DATA	=>	HPS_ENET_RX_DATA,
HPS_ENET_RX_DV	=>	HPS_ENET_RX_DV,
HPS_ENET_TX_DATA	=>	HPS_ENET_TX_DATA,
HPS_ENET_TX_EN	=>	HPS_ENET_TX_EN,
HPS_KEY	=>	HPS_KEY,
HPS_SD_CLK	=>	HPS_SD_CLK,
HPS_SD_CMD	=>	HPS_SD_CMD,
HPS_SD_DATA	=>	HPS_SD_DATA,
HPS_UART_RX	=>	HPS_UART_RX,
HPS_UART_TX	=>	HPS_UART_TX,
HPS_USB_CLKOUT	=>	HPS_USB_CLKOUT,
HPS_USB_DATA	=>	HPS_USB_DATA,
HPS_USB_DIR	=>	HPS_USB_DIR,
HPS_USB_NXT	=>	HPS_USB_NXT,
HPS_USB_STP	=>	HPS_USB_STP
        );

END MAIN;

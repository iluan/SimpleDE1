library IEEE;
use IEEE.STD_LOGIC_1164.all;
use ieee.numeric_std.all;

entity WRAP0 is
	port ( 
	--inserta aquí tus puertos
	);
end;
architecture synth of WRAP0 is
--inserta aquí tus señales y componentes
begin
--inserta aquí tus mapas de puerto, procesos y conexiones
end;
